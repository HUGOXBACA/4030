*********** LAB_2**************I
Is 0 1 4m
R0  1  2 12kohm
R1  2 0  12Kohms
R2  2 3 12Kohms
R3  1 3 12kohms
R4  3 0 12kohms


.TRAN 1m 5m
.PLOT  TRAN V(Is)
.PROBE
.END