****CSE4030Lab12****

Vs  1 0 PWL(0 0 0.1m 10) 
R1 1 2 1k
C1 2 0 10u

.TRAN 1ms 100ms
.PLOT TRAN V(1)
.PROBE 
.END