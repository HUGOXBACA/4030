****CSE4030Lab7pt2*****

Vs 0 1 DC 6V
R1 1 2  2k
R2 2 3  2k
R3 1 3 12k
R4 3 0 6k 



.Tran 1ms 7ms
.PLOT Tran V(1)
.PROBE
.END