******************Lab1_1**************************
Vs 1 0 9
R1 1 2 6
R2 2 0 3

.Tran 1m 5ms 
.PLOT Tran V(1)
.PROBE 
.END

