****CSE4030Lab10****

Vs 1 0 SIN(0 14.14 60 0 0 60) 
R1 1 2 2
L  2 0 5.3mH 

.Tran 2ms 100ms
.PLOT Tran V(1)
.PROBE
.END
