****CSE4030Lab11_pt2****

Vs 1 0 AC 0.01
E1 3 0 2 0 1000
C1 1 2 3.18nF
C2 4 0 79.58nF
R1 2 0 1000k
R2 3 4 100

.AC DEC 10 0.01 1000k 
.PLOT AC V(1)
.PROBE
.END 