*****test*****
Vs 1 0 DC 0.9mA
R1 1 2 60K
R2 2 0 40K
R3 20 80k

.Tran 1ms 5ms
.PLOT TRAN V(1) V(2)
.PROBE
.END