****CSE4030Lab13_pt1****

Vi 1 0 PWL(0 0 0.1m 1V )
R1 1 2 1
R2 2 0 1
L1 2 3  1
C1 3 0  4

.TRAN 1s 100s
.PLOT TRAN V(1)
.PROBE
.END
